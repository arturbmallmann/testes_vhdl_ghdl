package constantes is
	constant N : integer :=4;
end package;